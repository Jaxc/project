library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity IO_expander_APB is
  generic(
    pindex      : integer := 0;
    paddr       : integer := 0;
    pmask       : integer := 16#fff#
    );
  port (
    rstn  	: in  std_ulogic;
    clk   	: in  std_ulogic;
    apbi   	: in  apb_slv_in_type;
    apbo   	: out apb_slv_out_type;
    SDA		: inout STD_LOGIC;
    SCL_out	: out STD_LOGIC
  );                      
 
end entity IO_expander_APB;

architecture rtl of IO_expander_APB is

  -- APB related signals
  type adder_registers is record
    A       : std_logic_vector(31 downto 0);
    B       : std_logic_vector(31 downto 0);
    sum     : std_logic_vector(31 downto 0);
  end record;

  signal apb_reg    : adder_registers;
  signal apb_reg_in : adder_registers;
  
  signal A       : std_logic_vector(31 downto 0);
  signal B       : std_logic_vector(31 downto 0);
  signal sum     : std_logic_vector(31 downto 0);

	COMPONENT IO_explander_interface
	PORT(
		SCL : IN std_logic;
		rst : IN std_logic;
		I2C_slave_Address :in STD_LOGIC_VECTOR(6 downto 0);
		start_transmission : IN std_logic;
		Invector : IN std_logic_vector(7 downto 0);    
		SDA : INOUT std_logic;      
		IO_Ready : OUT std_logic;
		SCL_ena : OUT std_logic
		);
	END COMPONENT;

--constant REVISION       : amba_version_type := 0; 
constant pconfig        : apb_config_type := (
                        0 => ahb_device_reg ( VENDOR_OPENCORES, GAISLER_GPREG, 0, 0, 0),
                        1 => apb_iobar(paddr, pmask));

signal freq_cnt 	: integer range 0 to 499;
signal SCL 			: STD_LOGIC;

begin


	process(clk, rstn)
	begin
		if rstn = '0' then
			freq_cnt <= 0;
			SCL <= '0';
		elsif rising_edge(clk) then
			if freq_cnt = 499 then
				freq_cnt <= 0;
				SCL <= not (SCL);
			else
				freq_cnt <= freq_cnt + 1;
			end if;
		end if;
	end process;
SCL_out <= SCL;
	


	Inst_IO_explander_interface: IO_explander_interface PORT MAP(
		SCL => SCL,
		rst => rstn,
		I2C_slave_Address => "0000000",
		start_transmission => '1',
		IO_Ready => open,
		SCL_ena => open,
		Invector => "00000000",
		SDA => SDA
	);


end rtl;

